
module i_decode 
(

);

endmodule